module rcv_d(
        rcv_d_in1,
        rcv_d_in2,
        rcv_d_in3,
        rcv_d_out1,
        rcv_d_out2
        );
//---------------------------------------       
input        rcv_d_in1;
input        rcv_d_in2;
input        rcv_d_in3;   
output [7:0] rcv_d_out1; 
output       rcv_d_out2; 
//--------------------------------------- 
// synthesizable RTL code
always @(*)
   begin
       //-----
       //-----
   end
endmodule