module xmit_b(
        xmit_b_in1,
        xmit_b_in2,
        xmit_b_out1,
        xmit_b_out2      
        );
 
 //---------------------------------------       
 input [7:0]  xmit_b_in1;
 input        xmit_b_in2;
 output       xmit_b_out1;
 output       xmit_b_out2;
 //--------------------------------------- 
 // synthesizable RTL code
 always @(*)
    begin
        //-----
        //-----
    end
 
endmodule
